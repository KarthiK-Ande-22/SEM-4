module instr_mem(
    input [31:0] pc, 
    output reg [31:0] instr,
    input stall
);
    reg [31:0] memory [0:1023]; // 1K words of memory

    initial begin
        // memory[8]  = 32'b0000000_00011_00000_010_00100_0100011; // sd x3, 4(x0)
        // memory[9]  = 32'b0000000_00100_00000_010_00010_0000011; // ld x2, 4(x0)
        // memory[10] = 32'b0000000_00010_01001_000_00100_0110011; // add x4, x2, x9
        // memory[11] = 32'b0000000_00100_00110_000_00101_0110011; // add x5, x4, x6


        // memory[12]  = 32'b0000000_00010_00001_000_00001_0110011; // add x1, x1, x2
        // memory[13]  = 32'b0000000_00011_00001_000_00001_0110011; // add x1, x1, x3
        // memory[14] =  32'b0000000_00100_00001_000_00001_0110011; // add x1, x1, x4

        // memory[3] = 32'b0000000_00100_00110_000_00101_0110011; // add x5, x4, x6

        // memory[2] = 32'b0100000_00010_01001_000_01000_0110011; // sub x8, x2, x9 
        // memory[6] = 32'b0000000_01001_01101_110_01000_0110011; // or x8, x13, x9 
        // memory[5] = 32'b0000000_01000_00000_000_00001_0110011; // add x1, x0, x8   (Initialize x1 = 1)

        // branch checking

        // memory[1] = 32'b0000000_01001_01101_000_01001_0110011; // add x9, x13, x9
        // memory[0] = 32'b0000000_01000_00000_000_00001_0110011; // add x1, x0, x8   (Initialize x1 = 1)
        // memory[3] = 32'b0000000_00011_00011_000_01000_1100011; // beq x2, x3, loop (branching example) 
        // memory[4] = 32'b0000000_01001_01101_000_01001_0110011; // add x9, x13, x9 
        // memory[7] = 32'b0000000_01000_00000_000_00001_0110011; // add x1, x0, 4   (Initialize x1 = 1)
        // memory[2] = 32'b0000000_00100_00001_000_00001_0110011; // add x1, x7, x9
        
        // branch checking end 

        // memory[1] = 32'b0000000_00011_00001_000_00001_0110011; // add x9, x13, x9
        // memory[0] = 32'b0000000_00010_00001_000_00001_0110011; // add x1, x0, x8   (Initialize x1 = 1)

        memory[0] = 32'b0000000_00010_00100_000_00101_0110011; // add x5, x2, x4
        memory[1] = 32'b0000000_00101_00000_010_00100_0100011; // sd x5, 4(x0)
        memory[2] = 32'b0000000_00100_00000_010_00010_0000011; // ld x2, 4(x0)

        
    end

    always @(*) begin
        if(!stall)begin
            instr = memory[pc[6:0]>>2]; 
        end
        
    end
endmodule