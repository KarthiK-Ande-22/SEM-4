module instr_mem(
    input [31:0] pc, 
    output reg [31:0] instr,
    output reg [31:0] ifid_instr
);
    reg [31:0] memory [0:1023]; // 1K words of memory

    initial begin
        // memory[3] = 32'b0000000_00100_00000_000_00001_0110011; // addi x1, x0, 16   (Initialize x1 = 1)
        // memory[2] = 32'b0000000_10000_00000_000_00010_0010011; // addi x2, x0, 16  (Initialize x1 = 1)

        // memory[1] = 32'b0100000_01001_01101_000_01001_0110011; // sub x9, x13, x9
        // memory[0] = 32'b0000000_01001_01101_000_01001_0110011; // add x9, x13, x9  
        // memory[0]=32'b00000000000000010011001010000011; // ld x5, 0(x2)
        // memory[1]=32'b00000000000100010011001100000011;  // ld x6, 1(x2)
        // memory[2]=32'b00000000010100110000001000110011;  // add x4, x6, x5
        // memory[3]=32'b00000000001000010011001110000011; // ld x7, 2(x2)
        // memory[4]=32'b00000000011100100000001000110011;  // add x4, x4, x7
        // memory[5]=32'b00000000001100010011010000000011;  // ld x8, 3(x2)
        // memory[6]=32'b00000000100000100000001000110011;  // add x4, x4, x8
        // memory[7]=32'b00000000010000010011010010000011;  // ld x9, 4(x2)
        // memory[8]=32'b00000000100100100000001000110011;  // add x4, x4, x9
        // memory[9]=32'b00000000010000011011000000100011;  // sd x4, 0(x3)
        // memory[10]=32'b00000000000000011011010100000011;  // ld x10, 0(x3)
        // memory[11]=32'b00000000101001010000010100110011;  // add x10, x10, x10
        // memory[12]=32'b00000000101000011011000000100011;  // sd x10, 0(x3)
        // memory[0]  = 32'b0000000_00001_00000_000_00001_0010011; // addi x1, x0, 1   (Initialize x1 = 1)
        // memory[1]  = 32'b0000000_00001_00000_010_00001_0100011; // sd x1, 0(x0)     (Store Fib(1) = 1)
        // memory[2]  = 32'b0000000_00001_00010_000_00100_0110011; // add x4, x1, x2
        // memory[3]  = 32'b0100000_00011_01001_000_00101_0110011; // sub x5, x9, x3
        // memory[4]  = 32'b0000000_00100_00000_010_01000_0100011; // sd x4, 8(x0)
        // memory[5]  = 32'b0000000_00101_00000_010_10000_0100011; // sd x5, 16(x0)
        // memory[6]  = 32'b0000000_01001_00011_000_00100_0110011; // add x4, x9, x3
        // memory[7]  = 32'b0100000_00010_00001_000_00101_0110011; // sub x5, x1, x2
        // memory[8] = 32'b0000000_01000_00000_010_00100_0000011; // ld x4, 8(x0)
        // memory[9] = 32'b0000000_10000_00000_010_00101_0000011; // ld x5, 16(x0)
        // memory[10] = 32'b0000000_00101_00100_111_00110_0110011; // and x6, x4, x5
        // memory[11] = 32'b0000000_00101_00100_110_00111_0110011; // or x7, x4, x5
        // memory[12] = 32'b0000000_00101_00100_100_01000_0110011; // xor x8, x4, x5
        // memory[13]  = 32'b0000000_01111_00000_000_01101_0010011; // addi x13, x0, 15
        // memory[14]  = 32'b0000000_01111_00000_000_01110_0010011; // addi x14, x0, 15
        // memory[15] = 32'b0000000_01110_01110_000_10000_1100011; // beq x14, x14, loop (branching example)
        // memory[16] = 32'b0000000_01111_00000_000_01111_0010011; // addi x15, x0, 15
        // memory[17] = 32'b0000000_00010_00001_111_00110_0110011; // and x6, x1, x2
        // memory[18] = 32'b0000000_00010_00001_110_00111_0110011; // or x7, x1, x2
        // memory[19] = 32'b0000000_00010_00010_100_01000_0110011; // xor x8, x2, x2
        // memory[20] = 32'b00000000100000000011110000100011; // sd x8, 24(x0)
        // memory[21] = 32'b00000001100000000011010010000011; // ld x9, 24(x0)
        // memory[27] = 32'b0000000_11001_00000_010_01010_1111111; // exit

        $readmemb("general.txt", memory);
        $readmemb("general2.txt", memory);
        
        
    end

    always @(*) begin
        instr = memory[pc[6:0]>>2]; // Fetch instruction using word-aligned address
        ifid_instr = instr;
    end
endmodule