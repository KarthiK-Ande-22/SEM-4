module instr_mem(
    input [31:0] pc, 
    output reg [31:0] instr,
    input stall
);
    reg [31:0] memory [0:1023]; // 1K words of memory

    initial begin
        // memory[8]  = 32'b0000000_00011_00000_010_00100_0100011; // sd x3, 4(x0)
        // memory[9]  = 32'b0000000_00100_00000_010_00010_0000011; // ld x2, 4(x0)
        // memory[10] = 32'b0000000_00010_01001_000_00100_0110011; // add x4, x2, x9
        // memory[11] = 32'b0000000_00100_00110_000_00101_0110011; // add x5, x4, x6


        // memory[12]  = 32'b0000000_00010_00001_000_00001_0110011; // add x1, x1, x2
        // memory[13]  = 32'b0000000_00011_00001_000_00001_0110011; // add x1, x1, x3
        // memory[14] =  32'b0000000_00100_00001_000_00001_0110011; // add x1, x1, x4

        // memory[3] = 32'b0000000_00100_00110_000_00101_0110011; // add x5, x4, x6

        // memory[2] = 32'b0100000_00010_01001_000_01000_0110011; // sub x8, x2, x9 
        // memory[6] = 32'b0000000_01001_01101_110_01000_0110011; // or x8, x13, x9 
        // memory[5] = 32'b0000000_01000_00000_000_00001_0110011; // add x1, x0, x8   (Initialize x1 = 1)

        // branch checking

        // memory[1] = 32'b0000000_01001_01101_000_01001_0110011; // add x9, x13, x9
        // memory[0] = 32'b0000000_01000_00000_000_00001_0110011; // add x1, x0, x8   (Initialize x1 = 1)
        // memory[3] = 32'b0000000_00011_00011_000_01000_1100011; // beq x2, x3, loop (branching example) 
        // memory[4] = 32'b0000000_01001_01101_000_01001_0110011; // add x9, x13, x9 
        // memory[7] = 32'b0000000_01000_00000_000_00001_0110011; // add x1, x0, 4   (Initialize x1 = 1)
        // memory[2] = 32'b0000000_00100_00001_000_00001_0110011; // add x1, x7, x9
        
        // branch checking end 

        // memory[1] = 32'b0000000_00011_00001_000_00001_0110011; // add x9, x13, x9
        // memory[0] = 32'b0000000_00010_00001_000_00001_0110011; // add x1, x0, x8   (Initialize x1 = 1)

        // memory[0] = 32'b0000000_00010_00100_000_00101_0110011; // add x5, x2, x4
        // memory[1] = 32'b0000000_00101_00000_010_00100_0100011; // sd x5, 4(x0)
        // memory[2] = 32'b0000000_00100_00000_010_00010_0000011; // ld x2, 4(x0)

        // memory[0] = 32'b0000000_00010_00001_000_00001_0110011; // add x1, x1, x2
        // memory[1] = 32'b0000000_00011_00001_000_00001_0110011; // add x1, x1, x3
        // memory[2] = 32'b0000000_00100_00001_000_00001_0110011; // add x1, x1, x4
        // memory[7] = 32'b0000000_11001_00000_010_01010_1111111; // exit

        // memory[0]=32'b00000000000000010011001010000011; // ld x5, 0(x2)
        // memory[1]=32'b00000000000100010011001100000011;  // ld x6, 1(x2)
        // memory[2]=32'b00000000010100110000001000110011;  // add x4, x6, x5
        // memory[3]=32'b00000000001000010011001110000011; // ld x7, 2(x2)
        // memory[4]=32'b00000000011100100000001000110011;  // add x4, x4, x7
        // memory[5]=32'b00000000001100010011010000000011;  // ld x8, 3(x2)
        // memory[6]=32'b00000000100000100000001000110011;  // add x4, x4, x8
        // memory[7]=32'b00000000010000010011010010000011;  // ld x9, 4(x2)
        // memory[8]=32'b00000000100100100000001000110011;  // add x4, x4, x9
        // memory[9]=32'b00000000010000011011000000100011;  // sd x4, 0(x3)
        // memory[10]=32'b00000000000000011011010100000011;  // ld x10, 0(x3)
        // memory[11]=32'b00000000101001010000010100110011;  // add x10, x10, x10
        // memory[12]=32'b00000000101000011011000000100011;  // sd x10, 0(x3)
        // memory[17]=32'b00000000101000011011000001111111;  // sd x10, 0(x3)

        // memory[0]= 32'b0000000_00001_00000_000_00001_0010011;  //addi x1, x0, 1   (Initialize x1 = 1)
        // memory[1]= 32'b0000000_00001_00000_010_00001_0100011;  //sd x1, 0(x0)     (Store Fib(1) = 1)
        // memory[2]= 32'b0000000_00001_00000_000_00010_0010011;  //addi x2, x0, 1   (Initialize x2 = 1)
        // memory[3]= 32'b0000000_00010_00000_010_00010_0100011;  //sd x2, 8(x0)     (Store Fib(2) = 1)
        // memory[4]= 32'b0000000_00010_00000_000_00011_0010011;  //addi x3, x0, 2   (Counter x3 = 2)
        // memory[5]= 32'b0000000_01010_00000_000_01000_0010011;  //addi x8, x0, 10   (Loop limit N=6)
        // memory[6]= 32'b0000000_00001_00010_000_00100_0110011;  //add x4, x1, x2   (Fib(n) = x1 + x2)
        // memory[7]= 32'b0000000_00100_00000_010_00100_0100011;  //sd x4, 16(x0)    (Store Fib(n))
        // memory[8]= 32'b0000000_00010_00000_000_00001_0110011;  //add x1, x2, x0   (x1 = x2)
        // memory[9]= 32'b0000000_00100_00000_000_00010_0110011;  //add x2, x4, x0   (x2 = x4)
        // memory[10]= 32'b0000000_00001_00011_000_10100_0010011;  //addi x20, x3, 1   (Increment counter)
        // memory[11]= 32'b0000000_00000_10100_000_00011_0010011;  //addi x3, x20, 0   (Update counter)
        // memory[12]= 32'b0000000_00011_01000_000_00110_1100011;  //beq x3, x8, exit  (Exit if x3 == N)
        // memory[13]= 32'b1111111_00000_00000_000_10001_1100011;  //beq x0, x0, -32   (Jump back to loop)
        // memory[14]= 32'b0000000_00000_00000_000_00000_0000000;  //nop
        // memory[15]= 32'b0000000_00001_00000_000_01111_0010011;  //addi x15, x0, 1   (Final instruction)
        // memory[16]= 32'b0000000_00000_00000_000_00000_1111111;  //nop

        
        // memory[0]  = 32'b0000000_00001_00000_000_00001_0010011; // addi x1, x0, 1   (Initialize x1 = 1)
        // memory[1]  = 32'b0000000_00001_00000_010_00001_0100011; // sd x1, 0(x0)     (Store Fib(1) = 1)
        // memory[2]  = 32'b0000000_00001_00010_000_00100_0110011; // add x4, x1, x2
        // memory[3]  = 32'b0100000_00011_01001_000_00101_0110011; // sub x5, x9, x3
        // memory[4]  = 32'b0000000_00100_00000_010_01000_0100011; // sd x4, 8(x0)
        // memory[5]  = 32'b0000000_00101_00000_010_10000_0100011; // sd x5, 16(x0)
        // memory[6]  = 32'b0000000_01001_00011_000_00100_0110011; // add x4, x9, x3
        // memory[7]  = 32'b0100000_00010_00001_000_00101_0110011; // sub x5, x1, x2
        // memory[8] = 32'b0000000_01000_00000_010_00100_0000011; // ld x4, 8(x0)
        // memory[9] = 32'b0000000_10000_00000_010_00101_0000011; // ld x5, 16(x0)
        // memory[10] = 32'b0000000_00101_00100_111_00110_0110011; // and x6, x4, x5
        // memory[11] = 32'b0000000_00101_00100_110_00111_0110011; // or x7, x4, x5
        // memory[12] = 32'b0000000_00101_00100_100_01000_0110011; // xor x8, x4, x5
        // memory[13]  = 32'b0000000_01111_00000_000_01101_0010011; // addi x13, x0, 15
        // memory[14]  = 32'b0000000_01111_00000_000_01110_0010011; // addi x14, x0, 15
        // memory[15] = 32'b0000000_01110_01110_000_00100_1100011; // beq x13, x13, loop (branching example)
        // memory[16] = 32'b0000000_01110_00000_000_01111_0010011; // addi x15, x0, 14
        // memory[17] = 32'b0000000_00010_00001_111_00110_0110011; // and x6, x1, x2
        // memory[18] = 32'b0000000_00010_00001_110_00111_0110011; // or x7, x1, x2
        // memory[19] = 32'b0000000_00010_00010_100_01000_0110011; // xor x8, x2, x2
        // memory[20] = 32'b00000000100000000011110000100011; // sd x8, 24(x0)
        // memory[21] = 32'b00000001100000000011010010000011; // ld x9, 24(x0)
        // memory[27] = 32'b0000000_11001_00000_010_01010_1111111; // exit


        // $readmemb("hazard_fibbanocci.txt", memory);
        $readmemb("hazard_general1.txt", memory);
        // $readmemb("hazard_general2.txt", memory);
        // $readmemb("hazard_general3.txtt", memory);
        // $readmemb("hazard_double.txt", memory);

        
    end

    always @(*) begin
        if(!stall)begin
            instr = memory[pc[6:0]>>2]; 
        end
        
    end
endmodule